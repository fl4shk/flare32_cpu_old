`include "src/cpu_defines.svinc"


module Cpu(input wire clk,
	output a);


endmodule
