`include "src/misc_defines.svinc"
